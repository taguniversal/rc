module nash_permutation_tables (
    input wire [7:0] index,
    output reg [7:0] red_next_state,
    output reg red_transform,
    output reg [7:0] blue_next_state,
    output reg blue_transform
);

    always @* begin
        case (index)
            8'd0: begin red_next_state = 8'd63; red_transform = 1'b1; end
            8'd1: begin red_next_state = 8'd8; red_transform = 1'b1; end
            8'd2: begin red_next_state = 8'd52; red_transform = 1'b1; end
            8'd3: begin red_next_state = 8'd10; red_transform = 1'b0; end
            8'd4: begin red_next_state = 8'd118; red_transform = 1'b0; end
            8'd5: begin red_next_state = 8'd68; red_transform = 1'b1; end
            8'd6: begin red_next_state = 8'd93; red_transform = 1'b0; end
            8'd7: begin red_next_state = 8'd114; red_transform = 1'b0; end
            8'd8: begin red_next_state = 8'd54; red_transform = 1'b1; end
            8'd9: begin red_next_state = 8'd51; red_transform = 1'b0; end
            8'd10: begin red_next_state = 8'd3; red_transform = 1'b0; end
            8'd11: begin red_next_state = 8'd81; red_transform = 1'b0; end
            8'd12: begin red_next_state = 8'd37; red_transform = 1'b1; end
            8'd13: begin red_next_state = 8'd1; red_transform = 1'b0; end
            8'd14: begin red_next_state = 8'd21; red_transform = 1'b1; end
            8'd15: begin red_next_state = 8'd30; red_transform = 1'b0; end
            8'd16: begin red_next_state = 8'd92; red_transform = 1'b1; end
            8'd17: begin red_next_state = 8'd111; red_transform = 1'b1; end
            8'd18: begin red_next_state = 8'd35; red_transform = 1'b0; end
            8'd19: begin red_next_state = 8'd49; red_transform = 1'b0; end
            8'd20: begin red_next_state = 8'd79; red_transform = 1'b1; end
            8'd21: begin red_next_state = 8'd104; red_transform = 1'b1; end
            8'd22: begin red_next_state = 8'd24; red_transform = 1'b0; end
            8'd23: begin red_next_state = 8'd34; red_transform = 1'b1; end
            8'd24: begin red_next_state = 8'd5; red_transform = 1'b0; end
            8'd25: begin red_next_state = 8'd2; red_transform = 1'b0; end
            8'd26: begin red_next_state = 8'd38; red_transform = 1'b1; end
            8'd27: begin red_next_state = 8'd126; red_transform = 1'b0; end
            8'd28: begin red_next_state = 8'd121; red_transform = 1'b0; end
            8'd29: begin red_next_state = 8'd50; red_transform = 1'b1; end
            8'd30: begin red_next_state = 8'd7; red_transform = 1'b1; end
            8'd31: begin red_next_state = 8'd23; red_transform = 1'b1; end
            8'd32: begin red_next_state = 8'd46; red_transform = 1'b1; end
            8'd33: begin red_next_state = 8'd73; red_transform = 1'b1; end
            8'd34: begin red_next_state = 8'd42; red_transform = 1'b0; end
            8'd35: begin red_next_state = 8'd45; red_transform = 1'b0; end
            8'd36: begin red_next_state = 8'd83; red_transform = 1'b0; end
            8'd37: begin red_next_state = 8'd16; red_transform = 1'b0; end
            8'd38: begin red_next_state = 8'd120; red_transform = 1'b1; end
            8'd39: begin red_next_state = 8'd41; red_transform = 1'b0; end
            8'd40: begin red_next_state = 8'd95; red_transform = 1'b1; end
            8'd41: begin red_next_state = 8'd67; red_transform = 1'b0; end
            8'd42: begin red_next_state = 8'd60; red_transform = 1'b0; end
            8'd43: begin red_next_state = 8'd87; red_transform = 1'b1; end
            8'd44: begin red_next_state = 8'd85; red_transform = 1'b0; end
            8'd45: begin red_next_state = 8'd105; red_transform = 1'b1; end
            8'd46: begin red_next_state = 8'd70; red_transform = 1'b0; end
            8'd47: begin red_next_state = 8'd26; red_transform = 1'b1; end
            8'd48: begin red_next_state = 8'd117; red_transform = 1'b1; end
            8'd49: begin red_next_state = 8'd99; red_transform = 1'b1; end
            8'd50: begin red_next_state = 8'd80; red_transform = 1'b1; end
            8'd51: begin red_next_state = 8'd47; red_transform = 1'b1; end
            8'd52: begin red_next_state = 8'd77; red_transform = 1'b0; end
            8'd53: begin red_next_state = 8'd11; red_transform = 1'b1; end
            8'd54: begin red_next_state = 8'd29; red_transform = 1'b0; end
            8'd55: begin red_next_state = 8'd33; red_transform = 1'b1; end
            8'd56: begin red_next_state = 8'd43; red_transform = 1'b1; end
            8'd57: begin red_next_state = 8'd98; red_transform = 1'b0; end
            8'd58: begin red_next_state = 8'd103; red_transform = 1'b1; end
            8'd59: begin red_next_state = 8'd66; red_transform = 1'b0; end
            8'd60: begin red_next_state = 8'd6; red_transform = 1'b1; end
            8'd61: begin red_next_state = 8'd48; red_transform = 1'b1; end
            8'd62: begin red_next_state = 8'd78; red_transform = 1'b0; end
            8'd63: begin red_next_state = 8'd14; red_transform = 1'b1; end
            8'd64: begin red_next_state = 8'd96; red_transform = 1'b0; end
            8'd65: begin red_next_state = 8'd94; red_transform = 1'b0; end
            8'd66: begin red_next_state = 8'd127; red_transform = 1'b1; end
            8'd67: begin red_next_state = 8'd74; red_transform = 1'b1; end
            8'd68: begin red_next_state = 8'd28; red_transform = 1'b1; end
            8'd69: begin red_next_state = 8'd36; red_transform = 1'b1; end
            8'd70: begin red_next_state = 8'd123; red_transform = 1'b0; end
            8'd71: begin red_next_state = 8'd88; red_transform = 1'b1; end
            8'd72: begin red_next_state = 8'd76; red_transform = 1'b0; end
            8'd73: begin red_next_state = 8'd72; red_transform = 1'b0; end
            8'd74: begin red_next_state = 8'd62; red_transform = 1'b1; end
            8'd75: begin red_next_state = 8'd102; red_transform = 1'b0; end
            8'd76: begin red_next_state = 8'd53; red_transform = 1'b1; end
            8'd77: begin red_next_state = 8'd64; red_transform = 1'b0; end
            8'd78: begin red_next_state = 8'd69; red_transform = 1'b0; end
            8'd79: begin red_next_state = 8'd20; red_transform = 1'b1; end
            8'd80: begin red_next_state = 8'd71; red_transform = 1'b1; end
            8'd81: begin red_next_state = 8'd124; red_transform = 1'b1; end
            8'd82: begin red_next_state = 8'd31; red_transform = 1'b0; end
            8'd83: begin red_next_state = 8'd15; red_transform = 1'b1; end
            8'd84: begin red_next_state = 8'd86; red_transform = 1'b0; end
            8'd85: begin red_next_state = 8'd97; red_transform = 1'b0; end
            8'd86: begin red_next_state = 8'd116; red_transform = 1'b1; end
            8'd87: begin red_next_state = 8'd122; red_transform = 1'b1; end
            8'd88: begin red_next_state = 8'd82; red_transform = 1'b1; end
            8'd89: begin red_next_state = 8'd9; red_transform = 1'b0; end
            8'd90: begin red_next_state = 8'd32; red_transform = 1'b1; end
            8'd91: begin red_next_state = 8'd27; red_transform = 1'b1; end
            8'd92: begin red_next_state = 8'd106; red_transform = 1'b0; end
            8'd93: begin red_next_state = 8'd18; red_transform = 1'b1; end
            8'd94: begin red_next_state = 8'd56; red_transform = 1'b1; end
            8'd95: begin red_next_state = 8'd61; red_transform = 1'b1; end
            8'd96: begin red_next_state = 8'd110; red_transform = 1'b0; end
            8'd97: begin red_next_state = 8'd119; red_transform = 1'b1; end
            8'd98: begin red_next_state = 8'd57; red_transform = 1'b1; end
            8'd99: begin red_next_state = 8'd112; red_transform = 1'b0; end
            8'd100: begin red_next_state = 8'd100; red_transform = 1'b1; end
            8'd101: begin red_next_state = 8'd107; red_transform = 1'b1; end
            8'd102: begin red_next_state = 8'd65; red_transform = 1'b0; end
            8'd103: begin red_next_state = 8'd113; red_transform = 1'b1; end
            8'd104: begin red_next_state = 8'd19; red_transform = 1'b1; end
            8'd105: begin red_next_state = 8'd125; red_transform = 1'b1; end
            8'd106: begin red_next_state = 8'd91; red_transform = 1'b0; end
            8'd107: begin red_next_state = 8'd39; red_transform = 1'b1; end
            8'd108: begin red_next_state = 8'd55; red_transform = 1'b1; end
            8'd109: begin red_next_state = 8'd101; red_transform = 1'b0; end
            8'd110: begin red_next_state = 8'd75; red_transform = 1'b1; end
            8'd111: begin red_next_state = 8'd44; red_transform = 1'b1; end
            8'd112: begin red_next_state = 8'd115; red_transform = 1'b0; end
            8'd113: begin red_next_state = 8'd89; red_transform = 1'b1; end
            8'd114: begin red_next_state = 8'd109; red_transform = 1'b0; end
            8'd115: begin red_next_state = 8'd108; red_transform = 1'b0; end
            8'd116: begin red_next_state = 8'd22; red_transform = 1'b0; end
            8'd117: begin red_next_state = 8'd40; red_transform = 1'b0; end
            8'd118: begin red_next_state = 8'd90; red_transform = 1'b0; end
            8'd119: begin red_next_state = 8'd17; red_transform = 1'b1; end
            8'd120: begin red_next_state = 8'd0; red_transform = 1'b1; end
            8'd121: begin red_next_state = 8'd4; red_transform = 1'b1; end
            8'd122: begin red_next_state = 8'd13; red_transform = 1'b1; end
            8'd123: begin red_next_state = 8'd59; red_transform = 1'b1; end
            8'd124: begin red_next_state = 8'd12; red_transform = 1'b1; end
            8'd125: begin red_next_state = 8'd25; red_transform = 1'b1; end
            8'd126: begin red_next_state = 8'd58; red_transform = 1'b1; end
            8'd127: begin red_next_state = 8'd84; red_transform = 1'b1; end
            default: begin red_next_state = 8'd0; red_transform = 1'b0; end
        endcase
    end

    always @* begin
        case (index)
            8'd0: begin blue_next_state = 8'd30; blue_transform = 1'b1; end
            8'd1: begin blue_next_state = 8'd3; blue_transform = 1'b0; end
            8'd2: begin blue_next_state = 8'd112; blue_transform = 1'b1; end
            8'd3: begin blue_next_state = 8'd78; blue_transform = 1'b0; end
            8'd4: begin blue_next_state = 8'd20; blue_transform = 1'b1; end
            8'd5: begin blue_next_state = 8'd71; blue_transform = 1'b1; end
            8'd6: begin blue_next_state = 8'd54; blue_transform = 1'b1; end
            8'd7: begin blue_next_state = 8'd126; blue_transform = 1'b0; end
            8'd8: begin blue_next_state = 8'd17; blue_transform = 1'b0; end
            8'd9: begin blue_next_state = 8'd121; blue_transform = 1'b0; end
            8'd10: begin blue_next_state = 8'd107; blue_transform = 1'b0; end
            8'd11: begin blue_next_state = 8'd66; blue_transform = 1'b0; end
            8'd12: begin blue_next_state = 8'd86; blue_transform = 1'b1; end
            8'd13: begin blue_next_state = 8'd88; blue_transform = 1'b1; end
            8'd14: begin blue_next_state = 8'd9; blue_transform = 1'b0; end
            8'd15: begin blue_next_state = 8'd11; blue_transform = 1'b1; end
            8'd16: begin blue_next_state = 8'd45; blue_transform = 1'b1; end
            8'd17: begin blue_next_state = 8'd33; blue_transform = 1'b0; end
            8'd18: begin blue_next_state = 8'd4; blue_transform = 1'b1; end
            8'd19: begin blue_next_state = 8'd38; blue_transform = 1'b1; end
            8'd20: begin blue_next_state = 8'd91; blue_transform = 1'b1; end
            8'd21: begin blue_next_state = 8'd69; blue_transform = 1'b0; end
            8'd22: begin blue_next_state = 8'd35; blue_transform = 1'b0; end
            8'd23: begin blue_next_state = 8'd53; blue_transform = 1'b0; end
            8'd24: begin blue_next_state = 8'd109; blue_transform = 1'b0; end
            8'd25: begin blue_next_state = 8'd59; blue_transform = 1'b0; end
            8'd26: begin blue_next_state = 8'd28; blue_transform = 1'b0; end
            8'd27: begin blue_next_state = 8'd8; blue_transform = 1'b0; end
            8'd28: begin blue_next_state = 8'd123; blue_transform = 1'b0; end
            8'd29: begin blue_next_state = 8'd63; blue_transform = 1'b1; end
            8'd30: begin blue_next_state = 8'd10; blue_transform = 1'b0; end
            8'd31: begin blue_next_state = 8'd103; blue_transform = 1'b1; end
            8'd32: begin blue_next_state = 8'd29; blue_transform = 1'b1; end
            8'd33: begin blue_next_state = 8'd2; blue_transform = 1'b0; end
            8'd34: begin blue_next_state = 8'd22; blue_transform = 1'b1; end
            8'd35: begin blue_next_state = 8'd74; blue_transform = 1'b0; end
            8'd36: begin blue_next_state = 8'd58; blue_transform = 1'b1; end
            8'd37: begin blue_next_state = 8'd114; blue_transform = 1'b0; end
            8'd38: begin blue_next_state = 8'd76; blue_transform = 1'b1; end
            8'd39: begin blue_next_state = 8'd108; blue_transform = 1'b1; end
            8'd40: begin blue_next_state = 8'd125; blue_transform = 1'b0; end
            8'd41: begin blue_next_state = 8'd24; blue_transform = 1'b0; end
            8'd42: begin blue_next_state = 8'd51; blue_transform = 1'b0; end
            8'd43: begin blue_next_state = 8'd117; blue_transform = 1'b0; end
            8'd44: begin blue_next_state = 8'd49; blue_transform = 1'b0; end
            8'd45: begin blue_next_state = 8'd101; blue_transform = 1'b1; end
            8'd46: begin blue_next_state = 8'd18; blue_transform = 1'b1; end
            8'd47: begin blue_next_state = 8'd70; blue_transform = 1'b0; end
            8'd48: begin blue_next_state = 8'd21; blue_transform = 1'b1; end
            8'd49: begin blue_next_state = 8'd48; blue_transform = 1'b0; end
            8'd50: begin blue_next_state = 8'd110; blue_transform = 1'b0; end
            8'd51: begin blue_next_state = 8'd0; blue_transform = 1'b1; end
            8'd52: begin blue_next_state = 8'd116; blue_transform = 1'b1; end
            8'd53: begin blue_next_state = 8'd23; blue_transform = 1'b1; end
            8'd54: begin blue_next_state = 8'd104; blue_transform = 1'b1; end
            8'd55: begin blue_next_state = 8'd39; blue_transform = 1'b0; end
            8'd56: begin blue_next_state = 8'd40; blue_transform = 1'b1; end
            8'd57: begin blue_next_state = 8'd44; blue_transform = 1'b1; end
            8'd58: begin blue_next_state = 8'd94; blue_transform = 1'b1; end
            8'd59: begin blue_next_state = 8'd93; blue_transform = 1'b0; end
            8'd60: begin blue_next_state = 8'd1; blue_transform = 1'b1; end
            8'd61: begin blue_next_state = 8'd75; blue_transform = 1'b0; end
            8'd62: begin blue_next_state = 8'd127; blue_transform = 1'b0; end
            8'd63: begin blue_next_state = 8'd14; blue_transform = 1'b1; end
            8'd64: begin blue_next_state = 8'd32; blue_transform = 1'b0; end
            8'd65: begin blue_next_state = 8'd55; blue_transform = 1'b1; end
            8'd66: begin blue_next_state = 8'd52; blue_transform = 1'b1; end
            8'd67: begin blue_next_state = 8'd65; blue_transform = 1'b0; end
            8'd68: begin blue_next_state = 8'd99; blue_transform = 1'b0; end
            8'd69: begin blue_next_state = 8'd36; blue_transform = 1'b1; end
            8'd70: begin blue_next_state = 8'd50; blue_transform = 1'b0; end
            8'd71: begin blue_next_state = 8'd26; blue_transform = 1'b0; end
            8'd72: begin blue_next_state = 8'd111; blue_transform = 1'b1; end
            8'd73: begin blue_next_state = 8'd87; blue_transform = 1'b0; end
            8'd74: begin blue_next_state = 8'd27; blue_transform = 1'b0; end
            8'd75: begin blue_next_state = 8'd90; blue_transform = 1'b1; end
            8'd76: begin blue_next_state = 8'd62; blue_transform = 1'b0; end
            8'd77: begin blue_next_state = 8'd80; blue_transform = 1'b0; end
            8'd78: begin blue_next_state = 8'd13; blue_transform = 1'b1; end
            8'd79: begin blue_next_state = 8'd41; blue_transform = 1'b1; end
            8'd80: begin blue_next_state = 8'd6; blue_transform = 1'b1; end
            8'd81: begin blue_next_state = 8'd124; blue_transform = 1'b0; end
            8'd82: begin blue_next_state = 8'd84; blue_transform = 1'b0; end
            8'd83: begin blue_next_state = 8'd5; blue_transform = 1'b1; end
            8'd84: begin blue_next_state = 8'd92; blue_transform = 1'b1; end
            8'd85: begin blue_next_state = 8'd37; blue_transform = 1'b1; end
            8'd86: begin blue_next_state = 8'd15; blue_transform = 1'b1; end
            8'd87: begin blue_next_state = 8'd79; blue_transform = 1'b0; end
            8'd88: begin blue_next_state = 8'd64; blue_transform = 1'b0; end
            8'd89: begin blue_next_state = 8'd42; blue_transform = 1'b1; end
            8'd90: begin blue_next_state = 8'd96; blue_transform = 1'b0; end
            8'd91: begin blue_next_state = 8'd77; blue_transform = 1'b0; end
            8'd92: begin blue_next_state = 8'd12; blue_transform = 1'b1; end
            8'd93: begin blue_next_state = 8'd16; blue_transform = 1'b1; end
            8'd94: begin blue_next_state = 8'd7; blue_transform = 1'b1; end
            8'd95: begin blue_next_state = 8'd68; blue_transform = 1'b0; end
            8'd96: begin blue_next_state = 8'd46; blue_transform = 1'b0; end
            8'd97: begin blue_next_state = 8'd97; blue_transform = 1'b1; end
            8'd98: begin blue_next_state = 8'd102; blue_transform = 1'b1; end
            8'd99: begin blue_next_state = 8'd89; blue_transform = 1'b1; end
            8'd100: begin blue_next_state = 8'd106; blue_transform = 1'b0; end
            8'd101: begin blue_next_state = 8'd31; blue_transform = 1'b1; end
            8'd102: begin blue_next_state = 8'd119; blue_transform = 1'b0; end
            8'd103: begin blue_next_state = 8'd120; blue_transform = 1'b1; end
            8'd104: begin blue_next_state = 8'd47; blue_transform = 1'b0; end
            8'd105: begin blue_next_state = 8'd57; blue_transform = 1'b0; end
            8'd106: begin blue_next_state = 8'd60; blue_transform = 1'b1; end
            8'd107: begin blue_next_state = 8'd118; blue_transform = 1'b1; end
            8'd108: begin blue_next_state = 8'd83; blue_transform = 1'b1; end
            8'd109: begin blue_next_state = 8'd34; blue_transform = 1'b0; end
            8'd110: begin blue_next_state = 8'd98; blue_transform = 1'b0; end
            8'd111: begin blue_next_state = 8'd56; blue_transform = 1'b0; end
            8'd112: begin blue_next_state = 8'd105; blue_transform = 1'b0; end
            8'd113: begin blue_next_state = 8'd95; blue_transform = 1'b0; end
            8'd114: begin blue_next_state = 8'd43; blue_transform = 1'b1; end
            8'd115: begin blue_next_state = 8'd85; blue_transform = 1'b0; end
            8'd116: begin blue_next_state = 8'd122; blue_transform = 1'b0; end
            8'd117: begin blue_next_state = 8'd25; blue_transform = 1'b0; end
            8'd118: begin blue_next_state = 8'd67; blue_transform = 1'b1; end
            8'd119: begin blue_next_state = 8'd113; blue_transform = 1'b0; end
            8'd120: begin blue_next_state = 8'd81; blue_transform = 1'b1; end
            8'd121: begin blue_next_state = 8'd82; blue_transform = 1'b1; end
            8'd122: begin blue_next_state = 8'd115; blue_transform = 1'b1; end
            8'd123: begin blue_next_state = 8'd72; blue_transform = 1'b1; end
            8'd124: begin blue_next_state = 8'd100; blue_transform = 1'b1; end
            8'd125: begin blue_next_state = 8'd61; blue_transform = 1'b0; end
            8'd126: begin blue_next_state = 8'd19; blue_transform = 1'b1; end
            8'd127: begin blue_next_state = 8'd73; blue_transform = 1'b0; end
            default: begin blue_next_state = 8'd0; blue_transform = 1'b0; end
        endcase
    end
endmodule
